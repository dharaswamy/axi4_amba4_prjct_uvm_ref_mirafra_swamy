



//-------------------------------------------------------
//
//-------------------------------------------------------


//-------------------------------------------------------------------------------------------------------------------------------

// project : axi4 so: 
 `define AXI4_PROJECT 

// Project : axi3 :
// `define AXI3_PROJECT 

`define G_AXI_DATA_TYPE  bit 

//--------------------------------------------------------------------------------------------------
//   Write address channel signals widths : 
//--------------------------------------------------------------------------------------------------

//-------------------------------------------------------
//
//-------------------------------------------------------
   `define G_AXI_AWID_WIDTH  4
 
//-------------------------------------------------------
//
//-------------------------------------------------------
   `define G_AXI_AWADDR_WIDTH 32  // Default 
   
   //  `define G_AXI_AWADDR_WIDTH 64  // Default 

//-------------------------------------------------------
//
//-------------------------------------------------------
  `ifdef AXI3_PROJECT
  `define G_AXI_AWLEN_WIDTH 4
  `endif
  
  `ifdef AXI4_PROJECT
  `define G_AXI_AWLEN_WIDTH 8
  `endif

//-------------------------------------------------------
//
//-------------------------------------------------------
  `define G_AXI_AWSIZE_WIDTH 3 
  
//-------------------------------------------------------
//
//-------------------------------------------------------

  `define G_AXI_AWBURST_WIDTH 2
  
//-------------------------------------------------------
//
//-------------------------------------------------------

  `ifdef AXI3_PROJECT
  `define G_AXI_AWLOCK_WIDTH 2
   `endif

  `ifdef AXI4_PROJECT
     `define G_AXI_AWLOCK_WIDTH 1
    `endif
//-------------------------------------------------------
//
//-------------------------------------------------------
   `define G_AXI_AWCACHEE_WIDTH 4
//-------------------------------------------------------
//
//-------------------------------------------------------
  `define G_AXI_AWPROT_WIDTH 3
//-------------------------------------------------------
//
//-------------------------------------------------------
  `define G_AXI_AWQOS_WIDTH 4
//-------------------------------------------------------
//
//-------------------------------------------------------
  `define G_AXI_AWREGION_WIDTH 4

//-------------------------------------------------------

//-------------------------------------------------------

 `define G_AXI_AWUSER_WIDTH 1 

//--------------------------------------------------------------------------------------------------
//   Write DATA channel signals widths : 
//--------------------------------------------------------------------------------------------------

//-------------------------------------------------------
//
//-------------------------------------------------------
  `define  G_AXI_WID_WIDTH 4	

//-------------------------------------------------------
//
//-------------------------------------------------------

`define   G_AXI_WDATA_WIDTH 32 // Default

  // `define   G_AXI_WDATA_WIDTH 32 // Default
 //`define  G_AXI_WDATA_WIDTH 64 
 // `define  G_AXI_WDATA_WIDTH 128 
 //`define  G_AXI_WDATA_WIDTH 256
 //`define  G_AXI_WDATA_WIDTH 512
 //`define  G_AXI_WDATA_WIDTH 1024
 
//-------------------------------------------------------
//
//-------------------------------------------------------

 `define  G_AXI_WSTRB_WIDTH  `G_AXI_WDATA_WIDTH/8 


//-------------------------------------------------------
//
//-------------------------------------------------------
 `define G_AXI_WUSER_WIDTH 1
  
//--------------------------------------------------------------------------------------------------
//  Write response channel signals width : 
//--------------------------------------------------------------------------------------------------

//-------------------------------------------------------
//
//-------------------------------------------------------

 `define G_AXI_BID_WIDTH 4

//-------------------------------------------------------
//
//-------------------------------------------------------

`define G_AXI_BRESP_WIDTH 2

//-------------------------------------------------------
//
//-------------------------------------------------------

 `define G_AXI_BUSER_WIDTH 1

//--------------------------------------------------------------------------------------------------
//   Read address channel signals widths : 
//--------------------------------------------------------------------------------------------------

//-------------------------------------------------------
//
//-------------------------------------------------------
   `define G_AXI_ARID_WIDTH  4
 
//-------------------------------------------------------
//
//-------------------------------------------------------
   `define G_AXI_ARADDR_WIDTH 32  // Default 
   
   //  `define G_AXI_ARADDR_WIDTH 64  // Default 

//-------------------------------------------------------
//
//-------------------------------------------------------
  `ifdef AXI3_PROJECT
  `define G_AXI_ARLEN_WIDTH 4
  `endif

  `ifdef AXI4_PROJECT
  `define G_AXI_ARLEN_WIDTH 8
  `endif

//-------------------------------------------------------
//
//-------------------------------------------------------
  `define G_AXI_ARSIZE_WIDTH 3 
  
//-------------------------------------------------------
//
//-------------------------------------------------------

  `define G_AXI_ARBURST_WIDTH 2
  
//-------------------------------------------------------
//
//-------------------------------------------------------

  `ifdef AXI3_PROJECTl
  `define G_AXI_ARLOCK_WIDTH 2
  `endif

  `ifdef AXI4_PROJECT
  `define G_AXI_ARLOCK_WIDTH 1
   `endif

//-------------------------------------------------------
//
//-------------------------------------------------------
   `define G_AXI_ARCACHEE_WIDTH 4
//-------------------------------------------------------
//
//-------------------------------------------------------
  `define G_AXI_ARPROT_WIDTH 3
//-------------------------------------------------------
//
//-------------------------------------------------------
  `define G_AXI_ARQOS_WIDTH 4
//-------------------------------------------------------
//
//-------------------------------------------------------
  `define G_AXI_ARREGION_WIDTH 4

//-------------------------------------------------------
//
//-------------------------------------------------------
 `define G_AXI_ARUSER_WIDTH 1 

//--------------------------------------------------------------------------------------------------
//   Read DATA channel signals widths : 
//--------------------------------------------------------------------------------------------------

//-------------------------------------------------------
//
//-------------------------------------------------------
  `define  G_AXI_RID_WIDTH 4	

//-------------------------------------------------------
//
//-------------------------------------------------------
`define   G_AXI_RDATA_WIDTH 32 // Default

  // `define   G_AXI_RDATA_WIDTH 32 // Default
 //`define  G_AXI_RDATA_WIDTH 64 
 // `define  G_AXI_RDATA_WIDTH 128 
 //`define  G_AXI_RDATA_WIDTH 256
 //`define  G_AXI_RDATA_WIDTH 512
 //`define  G_AXI_RDATA_WIDTH 1024
 
//-------------------------------------------------------
//
//-------------------------------------------------------

`define G_AXI_RRESP_WIDTH 2
  
//-------------------------------------------------------
//
//-------------------------------------------------------
 `define G_AXI_RUSER_WIDTH 1


//================================================================================================================================



//-------------------------------------------------------
//
//-------------------------------------------------------




//-------------------------------------------------------
//
//-------------------------------------------------------




//-------------------------------------------------------
//
//-------------------------------------------------------

