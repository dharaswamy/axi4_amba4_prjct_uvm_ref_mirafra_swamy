

//--------------------------------------------------------------------------
//
//
//--------------------------------------------------------------------------




























//--------------------------------------------------------------------------
//
//
//--------------------------------------------------------------------------