
      
       

  //--------------------------------------------------------------------
  // Function/Task Name      : 
  // Parameters              :
  // Class  Name             :
  // Parent class Name       :
  // Usage or Purpose        :
  //--------------------------------------------------------------------
  
   //--------------------------------------------------------------------
  //
  //
  //
  //
  //--------------------------------------------------------------------
  

  //--------------------------------------------------------------------
  //
  //
  //
  //
  //--------------------------------------------------------------------
  

                             
                             